/****************************************************************************
 * wb_master_api_pkg.sv
 ****************************************************************************/

/**
 * Package: wb_master_api_pkg
 * 
 * TODO: Add package documentation
 */
package wb_master_api_pkg;
	
`ifdef HAVE_HDL_VIRTUAL_INTERFACE
	class wb_master_api;
		
		task reset();
			// TODO:
		endtask
		
		task response();
			// TODO:
		endtask
		
	endclass
`endif


endpackage


