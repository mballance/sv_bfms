
`include "uvm_macros.svh"

package wb_master_agent_pkg;
	import uvm_pkg::*;
	
	`include "wb_master_config.svh"
	`include "wb_master_seq_item.svh"
	`include "wb_master_driver.svh"
	`include "wb_master_monitor.svh"
	`include "wb_master_seq_base.svh"
	`include "wb_master_agent.svh"
endpackage



