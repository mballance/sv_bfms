/****************************************************************************
 * sv_bfms_utils_pkg.sv
 ****************************************************************************/

/**
 * Package: sv_bfms_utils_pkg
 * 
 * TODO: Add package documentation
 */
`include "uvm_macros.svh" 
package sv_bfms_utils_pkg;
	import uvm_pkg::*;
	import sv_bfms_api_pkg::*;
	
	`include "elf_loader.svh"

endpackage


