/****************************************************************************
 * wb_target_bfm.sv
 ****************************************************************************/
 
`ifndef WB_TARGET_BFM_NAME
`define WB_TARGET_BFM_NAME wb_target_bfm
`endif

/**
 * Interface: wb_target_bfm
 * 
 * TODO: Add interface documentation
 */
interface `WB_TARGET_BFM_NAME #(
		) ( );


endinterface


