/****************************************************************************
 * sv_bfms_api_dpi_pkg.sv
 ****************************************************************************/

/**
 * Package: sv_bfms_api_dpi_pkg
 * 
 * TODO: Add package documentation
 */
package sv_bfms_api_dpi_pkg;
	`include "sv_bfms_rw_api_dpi.svh"

endpackage


