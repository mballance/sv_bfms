/****************************************************************************
 * uart_serial_api_pkg.sv
 ****************************************************************************/

/**
 * Package: uart_serial_api_pkg
 * 
 * TODO: Add package documentation
 */
package uart_serial_api_pkg;
	
	class uart_serial_api;
		
	endclass


endpackage


